library verilog;
use verilog.vl_types.all;
entity cyclone_prim_dffe is
end cyclone_prim_dffe;
