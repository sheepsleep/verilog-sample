library verilog;
use verilog.vl_types.all;
entity sdr_tb is
end sdr_tb;
