module TFT_FullDisp(
input                     sys_clk  ,                //osc clock input
input                     sys_rst_n,                //ϵͳ��λ����

output  wire              LCD_SCL  ,                //LCDʹ���ź�
output  reg               LCD_SDA  ,                //LCD���������ߣ������ж���������Ϊ�����
output  reg               LCD_RS   ,                // PSB, 1 is  8 bit data mode
output  reg               LCD_CS   ,                // PSB, 1 is  8 bit data mode
output  reg               LCD_RST        
);   
