library verilog;
use verilog.vl_types.all;
entity TB_divide is
    generic(
        WIDTH           : integer := 10;
        SIZE            : integer := 8
    );
end TB_divide;
