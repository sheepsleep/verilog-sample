/**********************************************��Ȩ����*************************************************
**
**--------------------------------------------�ļ���Ϣ--------------------------------------------------
** �ļ����ƣ�        	74HC85.v
** ����޸����ڣ�    	2013-07-01
** ���°汾��        	V1.2
** ����������        	���һ��4λ�Ƚ����Ĺ���
**                                            
********************************************************************************************************/
module	compare4(
input	         [3:0]		key,				//	�Ƚ�ֵ
 
output  wire	[7:0]		LED 			   //	�ȽϽ�������
				);

// reg define
reg	[2:0]		f_out 			;
		
// wire define
wire	[4:0]		a_in  			;
wire	[3:0]		b_in  			;

//******************************************************************************
//  ģ�����ƣ�4λ�Ƚ���ģ��
//  �������������4λ�Ƚ����Ĺ���
//******************************************************************************
// assign  i_in is 3'b111 for run in our FPGA devlop board
assign i_in = 3'b111;                  //	��չ�����

assign a_in = { key[3:2], key[3:2] };  // ��һ��4λ�Ƚ�ֵ
assign b_in = { key[1:0], key[1:0] };  //	�ڶ���4λ�Ƚ�ֵ

assign LED = { 5'h0, f_out };          //	�ȽϽ��

// 74HC85 RTL Code
always@( * ) begin
	if ( a_in > b_in )
		 f_out =	3'b100;				   	//	���a����b			
	else if( a_in < b_in )
       f_out = 3'b010;					   //	���aС��b
	else begin
		case( i_in )
		3'b100:
				f_out = 3'b100;			   //	���a����b
		3'b010:
				f_out = 3'b010;			   //	���aС��b
		3'b001:						
				f_out = 3'b001;			   //	���a����b
  	   default:
				f_out = 3'b001; 		      //	���a����b
		endcase
	end
end

endmodule

// �Ա����̣�
// http://shop67541132.taobao.com
// http://shop69029874.taobao.com

