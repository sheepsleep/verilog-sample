/********************************��Ȩ����**************************************
**
**-------------------------------------------�ļ���Ϣ----------------------------------------------------------
** �ļ����ƣ�cmp.v
** ����������2λ�Ƚ���������
**           ���д��ڡ�С�ں͵��������жϹ���
** 
*******************************************************************************/
module cmp(
	A  ,				//�����ɿ��ؾ�����0�����£�1��δ����
	B  ,				//�����ɿ��ؾ�����0�����£�1��δ����
	F_M,				//���������0��������1��Ϩ��
	F_L,				//С�������0��������1��Ϩ��
	F_E					//���������0��������1��Ϩ��
	);						
input		[1:0]	A;		//����˿ڣ�2λ
input		[1:0]	B;		//����˿ڣ�2λ

output		F_M;			//����˿�
output		F_L;			//����˿�
output		F_E;			//����˿�

assign F_M = (A>B);			//ֱ�Ӹ�ֵ�����ڵ�ʱ������߼�1
assign F_L = (A<B);			//ֱ�Ӹ�ֵ��С�ڵ�ʱ������߼�1
assign F_E = (A==B);		//ֱ�Ӹ�ֵ�����ڵ�ʱ������߼�1

endmodule
