library verilog;
use verilog.vl_types.all;
entity tb_seg7 is
end tb_seg7;
