library verilog;
use verilog.vl_types.all;
entity print_task is
end print_task;
