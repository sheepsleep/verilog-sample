library verilog;
use verilog.vl_types.all;
entity tb_m4kram is
end tb_m4kram;
