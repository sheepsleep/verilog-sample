library verilog;
use verilog.vl_types.all;
entity SegLed_vlg_tst is
end SegLed_vlg_tst;
