library verilog;
use verilog.vl_types.all;
entity sld_signaltap is
    generic(
        sld_current_resource_width: integer := 0;
        sld_inversion_mask: string  := "0";
        sld_power_up_trigger: integer := 0;
        sld_advanced_trigger_6: string  := "NONE";
        sld_advanced_trigger_9: string  := "NONE";
        sld_advanced_trigger_7: string  := "NONE";
        sld_storage_qualifier_advanced_condition_entity: string  := "basic";
        sld_storage_qualifier_gap_record: integer := 0;
        sld_incremental_routing: integer := 0;
        sld_storage_qualifier_pipeline: integer := 0;
        sld_trigger_in_enabled: integer := 0;
        sld_state_bits  : integer := 5;
        sld_state_flow_use_generated: integer := 0;
        sld_inversion_mask_length: integer := 1;
        sld_data_bits   : integer := 1;
        sld_buffer_full_stop: integer := 1;
        sld_storage_qualifier_inversion_mask_length: integer := 0;
        sld_attribute_mem_mode: string  := "OFF";
        sld_storage_qualifier_mode: string  := "OFF";
        sld_state_flow_mgr_entity: string  := "state_flow_mgr_entity.vhd";
        sld_node_crc_loword: integer := 50132;
        sld_advanced_trigger_5: string  := "NONE";
        sld_trigger_bits: integer := 1;
        sld_storage_qualifier_bits: integer := 1;
        sld_advanced_trigger_10: string  := "NONE";
        sld_mem_address_bits: integer := 7;
        sld_advanced_trigger_entity: string  := "basic";
        sld_advanced_trigger_4: string  := "NONE";
        sld_trigger_level: integer := 10;
        sld_advanced_trigger_8: string  := "NONE";
        sld_ram_block_type: string  := "AUTO";
        sld_advanced_trigger_2: string  := "NONE";
        sld_advanced_trigger_1: string  := "NONE";
        sld_data_bit_cntr_bits: integer := 4;
        lpm_type        : string  := "sld_signaltap";
        sld_node_crc_bits: integer := 32;
        sld_sample_depth: integer := 16;
        sld_enable_advanced_trigger: integer := 0;
        sld_segment_size: integer := 0;
        sld_node_info   : integer := 0;
        sld_storage_qualifier_enable_advanced_condition: integer := 0;
        sld_node_crc_hiword: integer := 41394;
        sld_trigger_level_pipeline: integer := 1;
        sld_advanced_trigger_3: string  := "NONE";
        ela_status_bits : integer := 4;
        n_ela_instrs    : integer := 8
    );
    port(
        jtag_state_sdr  : in     vl_logic;
        ir_out          : out    vl_logic_vector;
        jtag_state_cdr  : in     vl_logic;
        ir_in           : in     vl_logic_vector;
        tdi             : in     vl_logic;
        acq_trigger_out : out    vl_logic_vector;
        jtag_state_uir  : in     vl_logic;
        acq_trigger_in  : in     vl_logic_vector;
        trigger_out     : out    vl_logic;
        storage_enable  : in     vl_logic;
        acq_data_out    : out    vl_logic_vector;
        acq_data_in     : in     vl_logic_vector;
        acq_storage_qualifier_in: in     vl_logic_vector;
        jtag_state_udr  : in     vl_logic;
        tdo             : out    vl_logic;
        clrn            : in     vl_logic;
        crc             : in     vl_logic_vector;
        jtag_state_e1dr : in     vl_logic;
        raw_tck         : in     vl_logic;
        usr1            : in     vl_logic;
        acq_clk         : in     vl_logic;
        shift           : in     vl_logic;
        ena             : in     vl_logic;
        trigger_in      : in     vl_logic;
        update          : in     vl_logic;
        rti             : in     vl_logic
    );
end sld_signaltap;
