library verilog;
use verilog.vl_types.all;
entity TB is
end TB;
