library verilog;
use verilog.vl_types.all;
entity altera_mf_hint_evaluation is
end altera_mf_hint_evaluation;
