library verilog;
use verilog.vl_types.all;
entity cyclone_and1 is
    port(
        y               : out    vl_logic;
        in1             : in     vl_logic
    );
end cyclone_and1;
