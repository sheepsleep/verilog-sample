library verilog;
use verilog.vl_types.all;
entity tb_sdrtest is
end tb_sdrtest;
