library verilog;
use verilog.vl_types.all;
entity altera_mf_memory_initialization is
end altera_mf_memory_initialization;
